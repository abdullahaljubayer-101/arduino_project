PK   �B�W�ӿ*  }J     cirkitFile.json͛�o�8������2ȡ���m���>�5���aP��H>Yn��/GV�8��3�n '��3����3�rt�m�E���'�m�	.��7�+���b��fٷˏ�Y���=쿬mX��붱M�L˸2�(�T&:����Mgƨ�(%�Z���j1�fuIS����G4uMS�i�	M=��gDl����D�$�<IDOٓD�$�>I�O"S�`l!MnC��<�T��<�y��J�Q��żɞc��HT���,��,V2,l�%�<u��pG��ᖈ=�"�@���{ bİ���)"����Sљ��u���WDt]u]ϸ7�r��е��zI�(�v�Mw�G���d��ĭ�þ:)�U����g1�L�پE
�`��X�D,V4����J�b%e���P�/��_�ï�X�,y�<K��bFR����y(���b�x(���b��Ŋ�b�C�bJ%x(V;��qB1�C��X�H�o��|�-`��3+Dj	V�%7����ȷD����oz�[j���mߙ1ݧ[+��J�bE�X�Y�$,VR+uL���+y�<�J�%��a�ð�X�P<S�x(���b�x(���b�C��X1�<+�Ŋ�b�"���>�ʋ�x���Z�N��V�ȥ�������/��sp�f�]���r�2�-��h��v����	e�3�3#��)=o����W��V��+��m?9
LSNq���X`��F�=���ȳ#�>� ,�+�u��i���VU�����K���%�NE�����5Q?&�'D����Q�!H%PR�T%BI�PR1�T%ġ��?@-�I���`L��	T0�
&P�*�@��J����Ȼ4�ġ$ru�~Q�TT0�3`zW�~�λ$b��ǃ����t��zW�'�ue��L]br��o0���(��S�Uñ)��RL�O�>�H2u���[Jl*����[Kl.��D��� Ԁ�6j j j j j j j j(�P�����P*�P��te��?�'�|����/<nwK��Wt�{���ۤ��!�H�ު��!9ŝ��9�K){p}�7�Vn�+$�����m����H��`^�f�Z�5e޺RyY7U�\՛W�t�I�*3Qa��:̫*m�dbc��([�n�^���Z�G-W���gL.���?Moܹ���e׮m��c>�o7u?�W�U�`�g�T�D����v�pyߺZ>(�J�M+����Q��2�R*7e��ԅ��4�N�+@͂���h�n0�0A7��+Vv��U"7B��b��X��њ$B<�H�EQ�ϊ�c���H+�>��']$��I�9���H��(>ד�����༖8�d�V}N��h}��x<��Q2��h�ϣh�ϣd�ϣh�ϣd�ϣd��;ɤ�Gє�Gф�Gɔ�Gє�Gє�Gф�w�)?��	?��?/������o˺���ߣ9�s�+�]7��k�黺���Dcn�;Jg�'�����{J�ŘSl����mnڻw�?���2��u�>ԛ:_�����o[w���])oM�uq��v�{n����~m�?��m�r�!�y�e&"�̥L��;�b0QlC�Wfn�	��6�8I*LZ��i��J�����$\�d���և�H���T���R�����Oo�r�:n&� ()�:�R�w;���:�'��������L@Xf����0��*��2�C��WJ�D����1�U<���|��w�mS�����E�/�!ep�!�Gn��q��e��i�J�C�rc�7���ȭ����#�X}��Ɩo���eg��ˇ������0�����������W=��ٵ��t�eݼ-�7��1۔Ϛ�,G[��{�96g�W��ۺ�/M3����0�}W]���p�m������~�Y���`6��������}�ag{����:xp8��{�������Ο�W̓�W��`���C�9r�V�y���V�.߽���r�d��s����O_���\a�N[1��wc�Ǡ��X4�^É�F�Պ�&8�j�������]���G�f�R�ߖ���Ҭ޴�o{{��	-��?PK   �B�W�ӿ*  }J             ��    cirkitFile.jsonPK      =   W    