PK   �wW�A��  i�     cirkitFile.json�][s���+)�+�5�z�ds�����lj� �X�̚udR��ֻq��I�æ�l"=��h4�ݍn �:��_�zYn�n���ޭ6����'���؇�����j��m��l������w����e����f�ֻ%%��tV�9ɸy�KQg�)���*]�e>����l�����Uu�q_!��W��J*m�K:�8t��2ôL}ˈ�W��\u���p�5���U'9�>A�G� �Gxd����<�+2n��t^��OA+��v����9�i$�	�	z�D=E��"QO)f�	��P�jgeP���0OQ��/VL���F��"�E�7�\o,�ތ+�Ȍ*t�)���*�+Ϋ�*�q���A-�<:U0���"Ld��¸�`��RU��lԗd\Yߊ��r�}e�TV��+i�Pu��Ĵ�3���:���T�UF+�|˥�l�lF�$e���%{�>�Z~�>ۼ$~�L��d�&3��3+m�\�+��&��Q}�#-�O�3*�o������d�K��s�#Hl��j�I��<�2Pl�4#���p�1�!u�=im�xŜ3��Cm�F+�B1�Ɍw��z�ب����@s�1��%F����Bj�ѺӲƴ�0-���)m�}�9RP�mT�1���cڎ)~��6J�خ��ƴ�2<$���d�m��o����	B���b�PC�Z!1}j9�� zGO} ��q�=Y��1u�| �`?�ߎ��rs��"���ﬨ�b���E	΋����;˛��O�E$�"�pQI��$\L.$OÆ�a��$~I�Ω�0lK�*V`ؤ�0I�a��$�i�4(�����]c�4(6��Ʈ��V	�Q���aR׵ðI�b��4�i�4(fgQ͈M+?hv+p�2�h�j�]IuijTX��TDhiZh6hZhf'pQU	rB�4�>YMe9��q���=���	I����4S��z�Dd5B��ӫH��D�q�i�B��������A��N¥��J���=�*e���G���/^N�2�8�/)N�2����LA}���^����t(��e@cj	�E�S��0ٴ,�hٴ)�F��.�)�u��;��b���nko�Q,<��K'�"�p�I��$\t.&��7zI��4�%i L� ���0I�a��$�i�D:8�i�4(�iPLӠ��A1M�b��,��Y��Xx.geG��\���bṜ���s9+8���rVp�%�,g�8���r���Xx.g8���r���X	P��i�{�#�G��I��9<�5���s9;��(����G��\�N58���rv��Q��os��o��I���mvE�|�e�uw��[�j�Z/7��mgW�ɯ��/a�a��H˘�=��H��Lo��y���3��J%�B&fi���x��>K�~3�2p��ٹ`Z���#-��cN����o��Ms��in��ȗ���k�D��f3�lPpL��	:���[�
���FG��-h:�C�;4�%X��R��'�m��I�z1\�뷨� z�i`�s �2fe?�� ~��Q�xTn��ͯ�Z�u5���2�ؾ�ch<&�sl�&x�]~���F����5R l��J  x���=
���@L�爝�G B��9b��@��'x��^ d�cR�g�u�A�y���$��xx�/V���� hȞn
��m� 5 Ԣ	�lڡ/!=������mo�7x���׺7 �W�7xqk��#�;z�#�ȼ�4=�� c��X���m�<�j�rD���6{�@l/2��`�)�" 3ۓ<G�/ 2����"A��<K�=$��_������d
/�ܯ*�8y���ȐJ1{vKD}��ϑ���D�W��Y� �7�lQ�����>mwM�%*��"V����X�,L	��S��i�MoV#� �a�?�s�#(68y`iP�cQL�(�XS,��l���l`���M�]��p�cq��O���E\g�70���������c��&��rTP���������݈t�@��� #v�:;�guz�0/�J�?�ӛ
PtZvf�7ٺ�^_ٻ��{d��yz�P�V�=2��=��Cȡ�~�'⛀��WD��_����U�Cp���v"�~ѧ7X�ށ����~ԧ7:���������ج�����Bp�<�/|�%h� �z��a���{X�ͺjtq�"5�Lw��k$ГP��4Ԡ�P�I��P��4Ԡ�5h��B�|m ��>��+@��N�Gک q; ~[�DG%�3�&di��� ��2�x�G���X���L������u�j���c6��S��ľ"�ε��@:�^�g8��:�4��{NQ!bL�u�c0
�/F�yG�������g��>��qG4�ྟ���p�����p���$�pۄ�:{ܑ��8(��~�`�M��Y�2n�`�7�iP_B�:�1��Yy��'yr����	�ro��.���O���JH[D�E�-��"��a�h�İH�ErX��"5,�m�����ȡ�d�gr�����i2�59����Ĭ�2>,;	�C��j����y�77�b�lUl�6<qQo�7��]@�E���3^*��.���MVH�ao�$�.%[��?����ǖ7��0GX~|3�������k������mw+�>߮��^ڻ�v����dm?��C�|����1-�ޯW��������ˏ�x������9_x�?��Vō;~�u��ںjv������l���-w�[��j�!�I��+[o�W�?�[W����	^���`���n��r�Yi4܄1'~>JIF��#�8��s����MVN��x5Q��^K����ܕyY��vv]�뀂���wp��{�f����r�-o\;��R�E������c�+����¡/_��V��v��j�����YP�O,8T����]H��a��9�f��\�v�@����kWeFXo��CC�cYj�j��Y^��
s��d@��߽�a��^T�����hA�5�\��� �3�Ȑ��S �; R��4~���j�s*��kGI�i[y0 ��Ԋe�z�˒g�Q�Q&��ynEM��l�d����n8&��q`:c��ɕ�G����?
�߫YoDn���^�$M}7��p����r>�֛�<S�|n�T���JM�R	�&�Q��j.�Xx���E
�!�1Ym�����Q�,@�����i� �����(Ct�>�AJ����0ϡ~���|,奡����}Slv���-��ω�}.�W'8�5���*WZ�lgBY�y��m������b����q J�l7>�Ý��K 1V��"g�*�y\s��(����˹"�[*j	� 5���~�f���Wo���uc�}oS� ��__Y��t�/��8��� ��<�&�*�{��rj�A���{�k�E�]惋�W��;�޻8��WL�"�}�t�jϋ�v�y��nh�b�H����z�r_��1�b��&����P��z���Q�@|����\P�(�����ד�S큜�,;�@S%jyV$�D^�̸��ڡ�m.��6Gz:� tv�xp[���0�0�u��@�}"�d�����.7!��'�ux����ꊱc]�D��t�Sj���?�r��Q(U��!M�����~�Ugh�lXN�9���-�^��p�ۂ�쵟&��;��C쵝36J�&��.?��~�S��������0~D��yS�~Onts��m�3l�p�ݍ��΍�[���Q��%g�#�f!S.�3Z�"��ֹ�K� t�
�`M����y���.��J�/奡��KH9l��U���6��@.$����,�"����w���r�+5���'׈>���䄅��oݚ�wx�S����?3�n��������xȤ|�0k�������;�w�B|��?x����j��j��$n��u5�
v��a��_~J)����t��nV��{�������ÇYH0�X�?5�.|zu��n@���G�3�*IA���{�9R����of�<�^0`�_
H�z��߂�Ɛj�j*˔���i�yR�AR ��Nf׿�R�BcSc@���;��R��@���}P��P�L�uʥ� v�:10Hw!0�A��)�ؙL����h�&?:E���;.�R��@���ө�)`�ƁQ��a����4Fj�S&��r>��8�:�){�'�J�����P�.`�0.��� �k0�T���뜚*%0�k>������@��qʃ��Z>Hr>���6�Χ�;S�
�9�Ȥ:G�� �d�R�D�g��߿tB@*�ʡ��Rȸ@���`��,��xhV�"%0xB��<��x4��k&�ѥ�|�Rts�@*��x)h�.ܾ2.����=��:�R�����:i^��S��άФZ���Bp�Π5���I��ڣRj�Td��_¨��t��@�8,Oct]�h	=Z�R-�K��w)�:g�@�R��p&�3�ʌ��;G�`DP�Y%ϓ�,�DSo�HZ/�>j��=�Y�ʃm@��w`�QuN����0�I]�IS�+ >C�f�l�%�]
���(̺Tz<u��n�D5:�`�AaV;�)a�@(�=/�d
�����m?�d�	?�b�L��2:Qo=�K��#&�QT���&�t���|���.�?�;��퓮��Q�TdB�Ӯt;�{,'�|�O�] ޥ�y�)4鵐n.	F5�k�9ɋ��0�� XH,]��������<joս`1b��cT�[j! ���zp�N�YQ�t{l*�.�] Z*�=*RԽ�Y�j|?-��D��r��|���

������=!�.s~A���Re��n��<�E{�Dt'S� �:<jDz�P�T�|O�zH0`�^�K� ��q�t�����F����ɉ0`T�KP'�`T{��kO����ٝۮ����* ��c�/W�ͮ��͟7��������f��PK   �wW�A��  i�             ��    cirkitFile.jsonPK      =       